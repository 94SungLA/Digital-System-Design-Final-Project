library verilog;
use verilog.vl_types.all;
entity alarm_clock_vlg_vec_tst is
end alarm_clock_vlg_vec_tst;
